module hello;
  $display("Hello github!");
endmodule
